// Depletion-mode n-type MOSFET

module dfet (x);

	inout x;

	pullup (x);

endmodule // dfet
